* C:\Users\Vlad\Desktop\Poli\ELTH\Lab2\Ex1\ex1.cir
V1 1 3 90
V2 4 3 50
V3 5 4 30
I1 1 0 6
R1 1 2 25
R2 0 3 12
R3 2 5 20
R4 3 2 10
R5 0 4 10
.dc V1 90 90 1
.print dc I(R1) I(R2) I(R3) I(R4) I(R5) V(I1)
.end

